// Actel Corporation Proprietary and Confidential
//  Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//  Revision Information:
// Jun09    Revision 4.1
// Aug10    Revision 4.2
// SVN Revision Information:
// SVN $Revision: 8508 $
// SVN $Date: 2009-06-15 16:49:49 -0700 (Mon, 15 Jun 2009) $
`define CUARTO  \
1 \
'b \
0
`define CUARTI  \
1 \
'b \
0
`define CUARTl  \
1 \
'b \
1
`define CUARTOI  \
1 \
'b \
1
`timescale 1ns/1ns
module
TOP_CoreUARTapb_0_Clock_gen
(
CUARTII
,
CUARTlI
,
CUARTOl
,
CUARTIl
,
CUARTll
,
BAUD_VAL_FRACTION
)
;
parameter
BAUD_VAL_FRCTN_EN
=
0
;
input
CUARTII
;
input
CUARTlI
;
input
[
12
:
0
]
CUARTOl
;
input
[
2
:
0
]
BAUD_VAL_FRACTION
;
output
CUARTIl
;
output
CUARTll
;
wire
CUARTIl
;
wire
CUARTll
;
reg
[
12
:
0
]
CUARTO0
;
reg
CUARTI0
;
reg
CUARTl0
;
reg
[
3
:
0
]
CUARTO1
;
generate
if
(
BAUD_VAL_FRCTN_EN
==
1
'b
1
)
begin
reg
CUARTI1
;
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
if
(
CUARTlI
==
1
'b
0
)
begin
CUARTI1
<=
1
'b
0
;
end
else
begin
if
(
CUARTO0
==
13
'b
0000000000001
)
begin
CUARTI1
<=
1
'b
1
;
end
else
begin
CUARTI1
<=
1
'b
0
;
end
end
end
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTl1
if
(
CUARTlI
===
1
'b
0
)
begin
CUARTO0
<=
13
'b
0000000000000
;
CUARTI0
<=
1
'b
0
;
end
else
begin
case
(
BAUD_VAL_FRACTION
)
3
'b
000
:
begin
if
(
CUARTO0
===
13
'b
0000000000000
)
begin
CUARTO0
<=
CUARTOl
;
CUARTI0
<=
1
'b
1
;
end
else
begin
CUARTO0
<=
CUARTO0
-
1
'b
1
;
CUARTI0
<=
1
'b
0
;
end
end
3
'b
001
:
begin
if
(
CUARTO0
==
13
'b
0000000000000
)
begin
if
(
(
CUARTO1
[
2
:
0
]
==
3
'b
111
)
&&
(
CUARTI1
==
1
'b
1
)
)
begin
CUARTO0
<=
CUARTO0
;
CUARTI0
<=
1
'b
0
;
end
else
begin
CUARTO0
<=
CUARTOl
;
CUARTI0
<=
1
'b
1
;
end
end
else
begin
CUARTO0
<=
CUARTO0
-
1
'b
1
;
CUARTI0
<=
1
'b
0
;
end
end
3
'b
010
:
begin
if
(
CUARTO0
==
13
'b
0000000000000
)
begin
if
(
(
CUARTO1
[
1
:
0
]
==
2
'b
11
)
&&
(
CUARTI1
==
1
'b
1
)
)
begin
CUARTO0
<=
CUARTO0
;
CUARTI0
<=
1
'b
0
;
end
else
begin
CUARTO0
<=
CUARTOl
;
CUARTI0
<=
1
'b
1
;
end
end
else
begin
CUARTO0
<=
CUARTO0
-
1
'b
1
;
CUARTI0
<=
1
'b
0
;
end
end
3
'b
011
:
begin
if
(
CUARTO0
==
13
'b
0000000000000
)
begin
if
(
(
(
(
CUARTO1
[
2
]
==
1
'b
1
)
||
(
CUARTO1
[
1
]
==
1
'b
1
)
)
&&
(
CUARTO1
[
0
]
==
1
'b
1
)
)
&&
(
CUARTI1
==
1
'b
1
)
)
begin
CUARTO0
<=
CUARTO0
;
CUARTI0
<=
1
'b
0
;
end
else
begin
CUARTO0
<=
CUARTOl
;
CUARTI0
<=
1
'b
1
;
end
end
else
begin
CUARTO0
<=
CUARTO0
-
1
'b
1
;
CUARTI0
<=
1
'b
0
;
end
end
3
'b
100
:
begin
if
(
CUARTO0
==
13
'b
0000000000000
)
begin
if
(
(
CUARTO1
[
0
]
==
1
'b
1
)
&&
(
CUARTI1
==
1
'b
1
)
)
begin
CUARTO0
<=
CUARTO0
;
CUARTI0
<=
1
'b
0
;
end
else
begin
CUARTO0
<=
CUARTOl
;
CUARTI0
<=
1
'b
1
;
end
end
else
begin
CUARTO0
<=
CUARTO0
-
1
'b
1
;
CUARTI0
<=
1
'b
0
;
end
end
3
'b
101
:
begin
if
(
CUARTO0
==
13
'b
0000000000000
)
begin
if
(
(
(
(
CUARTO1
[
2
]
==
1
'b
1
)
&&
(
CUARTO1
[
1
]
==
1
'b
1
)
)
||
(
CUARTO1
[
0
]
==
1
'b
1
)
)
&&
(
CUARTI1
==
1
'b
1
)
)
begin
CUARTO0
<=
CUARTO0
;
CUARTI0
<=
1
'b
0
;
end
else
begin
CUARTO0
<=
CUARTOl
;
CUARTI0
<=
1
'b
1
;
end
end
else
begin
CUARTO0
<=
CUARTO0
-
1
'b
1
;
CUARTI0
<=
1
'b
0
;
end
end
3
'b
110
:
begin
if
(
CUARTO0
==
13
'b
0000000000000
)
begin
if
(
(
(
CUARTO1
[
1
]
==
1
'b
1
)
||
(
CUARTO1
[
0
]
==
1
'b
1
)
)
&&
(
CUARTI1
==
1
'b
1
)
)
begin
CUARTO0
<=
CUARTO0
;
CUARTI0
<=
1
'b
0
;
end
else
begin
CUARTO0
<=
CUARTOl
;
CUARTI0
<=
1
'b
1
;
end
end
else
begin
CUARTO0
<=
CUARTO0
-
1
'b
1
;
CUARTI0
<=
1
'b
0
;
end
end
3
'b
111
:
begin
if
(
CUARTO0
==
13
'b
0000000000000
)
begin
if
(
(
(
(
CUARTO1
[
1
]
==
1
'b
1
)
||
(
CUARTO1
[
0
]
==
1
'b
1
)
)
||
(
CUARTO1
[
2
:
0
]
==
3
'b
100
)
)
&&
(
CUARTI1
==
1
'b
1
)
)
begin
CUARTO0
<=
CUARTO0
;
CUARTI0
<=
1
'b
0
;
end
else
begin
CUARTO0
<=
CUARTOl
;
CUARTI0
<=
1
'b
1
;
end
end
else
begin
CUARTO0
<=
CUARTO0
-
1
'b
1
;
CUARTI0
<=
1
'b
0
;
end
end
default
:
begin
if
(
CUARTO0
===
13
'b
0000000000000
)
begin
CUARTO0
<=
CUARTOl
;
CUARTI0
<=
1
'b
1
;
end
else
begin
CUARTO0
<=
CUARTO0
-
1
'b
1
;
CUARTI0
<=
1
'b
0
;
end
end
endcase
end
end
end
else
if
(
BAUD_VAL_FRCTN_EN
==
1
'b
0
)
begin
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTl1
if
(
CUARTlI
===
1
'b
0
)
begin
CUARTO0
<=
13
'b
0000000000000
;
CUARTI0
<=
1
'b
0
;
end
else
begin
if
(
CUARTO0
===
13
'b
0000000000000
)
begin
CUARTO0
<=
CUARTOl
;
CUARTI0
<=
1
'b
1
;
end
else
begin
CUARTO0
<=
CUARTO0
-
1
'b
1
;
CUARTI0
<=
1
'b
0
;
end
end
end
end
endgenerate
always
@
(
posedge
CUARTII
or
negedge
CUARTlI
)
begin
:
CUARTOOI
if
(
CUARTlI
===
1
'b
0
)
begin
CUARTO1
<=
4
'b
0000
;
CUARTl0
<=
1
'b
0
;
end
else
begin
if
(
CUARTI0
===
1
'b
1
)
begin
CUARTO1
<=
CUARTO1
+
1
'b
1
;
if
(
CUARTO1
===
4
'b
1111
)
begin
CUARTl0
<=
1
'b
1
;
end
else
begin
CUARTl0
<=
1
'b
0
;
end
end
end
end
assign
CUARTll
=
CUARTl0
&
CUARTI0
;
assign
CUARTIl
=
CUARTI0
;
endmodule
